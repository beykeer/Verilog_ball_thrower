module Ball_thrower()






endmodule 