module ball(clk, rst, update, xlength, ylength, ball);



endmodule 