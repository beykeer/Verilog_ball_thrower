module field_generate()













endmodule 